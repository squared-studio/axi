// Description here
// Author : name (email)
// This file is part of squared-studio:axi
// Copyright (c) 2025 squared-studio
// Licensed under the MIT License
// See LICENSE file in the project root for full license information

`include "axi4l_typedef.svh"
`include "vip/axi4l_pkg.sv"
`include "vip/axi4l_pkg_macros.svh"

module axi4l_pkg_tb;

  `define ENABLE_DUMPFILE

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "vip/tb_ess.sv"

  // AXI4L VIP CLASSES IMPORT
  `IMPORT_AXI4L_PKG_CLASSES

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  `AXI4L_T(main, 32, 64)

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // generates static task start_clk_i with tHigh:4ns tLow:6ns
  `CREATE_CLK(clk_i, 5ns, 5ns)

  logic arst_ni = 1;

  main_req_t req;
  main_resp_t resp;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INTERFACES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  `AXI4L_VIP(man, 1, clk_i, arst_ni, req, resp)
  `AXI4L_VIP(sub, 0, clk_i, arst_ni, req, resp)

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-CLASSES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  task static apply_reset();
    #100;
    arst_ni <= 0;
    #100;
    arst_ni <= 1;
    #100;
  endtask

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin  // main initial

    apply_reset();
    start_clk_i();

    sub_dvr.failure_odds = 10;

    man_dvr.start();
    sub_dvr.start();
    man_mon.start();

    @ (posedge clk_i);

    repeat (10) begin
      man_seq_item_t item;
      item = new();
      item.randomize();
      item._type = 1;
      // $display("\n%s\n", item.to_string());
      man_dvr_mbx.put(item);
      repeat (1) @(posedge clk_i);
      item = new item;
      item._type = 0;
      // $display("\n%s\n", item.to_string());
      man_dvr_mbx.put(item);
    end

    fork
      man_mon.wait_cooldown();
      sub_mon.wait_cooldown();
    join

    while (man_mon_mbx.num()) begin
      man_resp_item_t item;
      man_mon_mbx.get(item);
      $display("\n%s\n", item.to_string());
    end

    $finish;

  end

endmodule
