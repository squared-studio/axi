/*
Write a markdown documentation for this systemverilog module:
Author : Foez Ahmed (foez.official@gmail.com)
*/

`include "axi_grid_interfacing.svh"

module axi_grid_mni #(
    parameter type      req_t          = axi_default_param_pkg::mni_req_t,
    parameter type      resp_t         = axi_default_param_pkg::mni_resp_t,
    parameter type      grid_id_t      = axi_default_param_pkg::grid_id_t,
    parameter type      grid_aw_chan_t = axi_default_param_pkg::grid_aw_chan_t,
    parameter type      grid_w_chan_t  = axi_default_param_pkg::grid_w_chan_t,
    parameter type      grid_b_chan_t  = axi_default_param_pkg::grid_b_chan_t,
    parameter type      grid_ar_chan_t = axi_default_param_pkg::grid_ar_chan_t,
    parameter type      grid_r_chan_t  = axi_default_param_pkg::grid_r_chan_t,
    parameter grid_id_t NI_ID          = 0
) (
    input  logic  clk_i,
    input  logic  arst_ni,
    output req_t  req_o,
    input  resp_t resp_i,
    `AXI_GRID_MODULE_PORTS
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS GENERATED
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INITIAL CHECKS
  //////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef SIMULATION
`endif  // SIMULATION

endmodule
