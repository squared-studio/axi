/*
Write a markdown documentation for this systemverilog module:
Author : Foez Ahmed (foez.official@gmail.com)
*/

`include "axi_default_param_pkg.sv"

module axi_grid_vh_join #(
    parameter type      grid_id_t = axi_default_param_pkg::grid_id_t,
    parameter type      chan_t    = axi_default_param_pkg::grid_id_t,
    parameter grid_id_t NI_ID     = 0
) (
    input logic clk_i,
    input logic arst_ni,

    input  grid_id_t v_did_i,
    input  grid_id_t v_sid_i,
    input  chan_t    v_chan_i,
    input  logic     v_valid_i,
    output logic     v_ready_o,

    input  grid_id_t h_did_i,
    input  grid_id_t h_sid_i,
    input  chan_t    h_chan_i,
    input  logic     h_valid_i,
    output logic     h_ready_o,

    output grid_id_t did_o,
    output grid_id_t sid_o,
    output chan_t    chan_o,
    output logic     valid_o,
    input  logic     ready_i
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS GENERATED
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INITIAL CHECKS
  //////////////////////////////////////////////////////////////////////////////////////////////////

endmodule
